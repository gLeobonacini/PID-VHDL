Conversor_Int_Float_inst : Conversor_Int_Float PORT MAP (
		aclr	 => aclr_sig,
		clock	 => clock_sig,
		dataa	 => dataa_sig,
		result	 => result_sig
	);
